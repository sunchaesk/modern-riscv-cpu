
module riscv (

              );


endmodule
